--
--library IEEE;
--use IEEE.STD_LOGIC_1164.all;
-- 
--entity demux_1to4 is
-- port(
-- 
-- F : in STD_LOGIC;
-- S0,S1: in STD_LOGIC;
-- A,B,C,D: out STD_LOGIC
-- );
--end demux_1to4;
-- 
--architecture bhv of demux_1to4 is
--begin
--process (F,S0,S1) is
--begin
-- if (S0 ='0' and S1 = '0') then
-- A <= F;
-- elsif (S0 ='1' and S1 = '0') then
-- B <= F;
-- elsif (S0 ='0' and S1 = '1') then
-- C <= F;
-- else
-- D <= F;
-- end if;
-- 
--end process;
--end bhv;
library IEEE;

use IEEE.STD_LOGIC_1164.ALL;

use IEEE.STD_LOGIC_ARITH.ALL;

use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity DEMUX is

Port ( I : in  STD_LOGIC_vector(7 downto 0);

S : in STD_LOGIC_VECTOR (1 downto 0);

Y : out STD_LOGIC_VECTOR (31 downto 0));

end DEMUX;

architecture Behavioral of DEMUX is

begin

process (I, S)

begin

if (S <= "00") then

Y(7 downto 0)<=I ;

elsif (S <= "01") then

Y(15 downto 8) <= I ;

elsif (S <= "10") then

Y(23 downto 16) <= I ;

else

Y(31 downto 24) <= I ;

end if;

end process;

end Behavioral;